module registerFile(
	input [63:0] data,
	input [4:0] rs1,rs2,rd,
	input regWrite, clk, reset,
	output reg [63:0] readData1, readData2
);

reg [63:0] registers [31:0];

initial
begin
	registers[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	registers[1] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
	registers[2] = 64'b0000000000000000000000000000000000000000000000000000000000000010;
	registers[3] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
	registers[4] = 64'b0000000000000000000000000000000000000000000000000000000000000100;
	registers[5] = 64'b0000000000000000000000000000000000000000000000000000000000000101;
	registers[6] = 64'b0000000000000000000000000000000000000000000000000000000000000110;
	registers[7] = 64'b0000000000000000000000000000000000000000000000000000000000000111;
	registers[8] = 64'b0000000000000000000000000000000000000000000000000000000000001000;
	registers[9] = 64'b0000000000000000000000000000000000000000000000000000000000001001;
	registers[10] = 64'b0000000000000000000000000000000000000000000000000000000000001010;
	registers[11] = 64'b0000000000000000000000000000000000000000000000000000000000001011;
	registers[12] = 64'b0000000000000000000000000000000000000000000000000000000000001100;
	registers[13] = 64'b0000000000000000000000000000000000000000000000000000000000001101;
	registers[14] = 64'b0000000000000000000000000000000000000000000000000000000000001110;
	registers[15] = 64'b0000000000000000000000000000000000000000000000000000000000001111;
	registers[16] = 64'b0000000000000000000000000000000000000000000000000000000000010000;
	registers[17] = 64'b0000000000000000000000000000000000000000000000000000000000010001;
	registers[18] = 64'b0000000000000000000000000000000000000000000000000000000000010010;
	registers[19] = 64'b0000000000000000000000000000000000000000000000000000000000010011;
	registers[20] = 64'b0000000000000000000000000000000000000000000000000000000000010100;
	registers[21] = 64'b0000000000000000000000000000000000000000000000000000000000010101;
	registers[22] = 64'b0000000000000000000000000000000000000000000000000000000000010110;
	registers[23] = 64'b0000000000000000000000000000000000000000000000000000000000010111;
	registers[24] = 64'b0000000000000000000000000000000000000000000000000000000000011000;
	registers[25] = 64'b0000000000000000000000000000000000000000000000000000000000011001;
	registers[26] = 64'b0000000000000000000000000000000000000000000000000000000000011010;
	registers[27] = 64'b0000000000000000000000000000000000000000000000000000000000011011;
	registers[28] = 64'b0000000000000000000000000000000000000000000000000000000000011100;
	registers[29] = 64'b0000000000000000000000000000000000000000000000000000000000011101;
	registers[30] = 64'b0000000000000000000000000000000000000000000000000000000000011110;
	registers[31] = 64'b0000000000000000000000000000000000000000000000000000000000011111;
end


//Writing data operation:
always @ (posedge clk)
begin 
	registers[rd] <= data;
end

//Reading data operation: 
always @ (negedge clk)
begin 
	if (reset)
	begin
		readData1 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
		readData2 = 64'b0000000000000000000000000000000000000000000000000000000000000000;	
	end
	else
	begin
		readData1 <= registers[rs1];
		readData2 <= registers[rs2];
	end
end
endmodule